package CPUpack;

endpackage